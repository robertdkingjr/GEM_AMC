----------------------------------------------------------------------------------
-- Company: TAMU, a lot of this is taken from WU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date: 04/24/2016 04:52:35 AM
-- Module Name: TTC
-- Project Name: GEM_AMC
-- Description: Locks to TTC clock and decodes TTC commands from the backplane link. Also provides various controls and counters to be used for configuration, diagnostics and daq   
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

library UNISIM;
use UNISIM.VComponents.all;

use work.ctp7_utils_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.gem_pkg.all;
use work.synchronizer.all;
use work.ttc_clocks.all;
use work.ttc_cmd.all;
use work.ipbus_slave.all;
use work.ipb_addr_decode.all;
use work.registers.all;

--============================================================================
--                                                          Entity declaration
--============================================================================

entity ttc is
    port(
        -- reset
        reset_i           : in  std_logic;

        -- TTC backplane clock and data signals
        clk_40_ttc_p_i    : in  std_logic;
        clk_40_ttc_n_i    : in  std_logic;
        ttc_data_p_i      : in  std_logic;
        ttc_data_n_i      : in  std_logic;

        -- TTC clocks (40, 80, 160, 240, 320)
        ttc_clks_o        : out t_ttc_clks;

        -- TTC commands
        ttc_cmds_o        : out t_ttc_cmds;
    
        -- DAQ counters (L1A ID, Orbit ID, BX ID)
        ttc_daq_cntrs_o   : out t_ttc_daq_cntrs;

        -- IPbus
        ipb_reset_i       : in  std_logic;
        ipb_clk_i         : in  std_logic;
        ipb_mosi_i        : in  ipb_wbus;
        ipb_miso_o        : out ipb_rbus
    );

end ttc;

--============================================================================
--                                                        Architecture section
--============================================================================
architecture ttc_arch of ttc is

    --============================================================================
    --                                                         Signal declarations
    --============================================================================

    signal reset        : std_logic;
    signal reset_local  : std_logic;

    -- clocks
    signal clk_40  : std_logic;
    signal clk_80  : std_logic;
    signal clk_160 : std_logic;
    signal clk_240 : std_logic;
    signal clk_320 : std_logic;

    -- commands
    signal ttc_cmd : std_logic_vector(7 downto 0);
    signal ttc_l1a : std_logic;

    signal l1a_cmd        : std_logic;
    signal bc0_cmd        : std_logic;
    signal ec0_cmd        : std_logic;
    signal resync_cmd     : std_logic;
    signal oc0_cmd        : std_logic;
    signal start_cmd      : std_logic;
    signal stop_cmd       : std_logic;
    signal hard_reset_cmd : std_logic;
    signal calpulse_cmd   : std_logic;
    signal test_sync_cmd  : std_logic;

    -- daq counters
    signal l1id_cnt  : std_logic_vector(23 downto 0);
    signal orbit_cnt : std_logic_vector(15 downto 0);
    signal bx_cnt    : std_logic_vector(11 downto 0);

    -- control and status
    signal ttc_ctrl         : t_ttc_ctrl;
    signal ttc_status       : t_ttc_status;    

    -- stats
    constant C_NUM_OF_DECODED_TTC_CMDS : integer := 10;
    signal ttc_cmds_arr              : std_logic_vector(C_NUM_OF_DECODED_TTC_CMDS - 1 downto 0);
    signal ttc_cmds_cnt_arr          : t_slv_arr_32(C_NUM_OF_DECODED_TTC_CMDS - 1 downto 0);

    -- ttc mini spy
    signal ttc_spy_buffer    : std_logic_vector(31 downto 0) := (others => '1');
    signal ttc_spy_pointer   : integer range 0 to 31         := 0;
    signal ttc_spy_reset     : std_logic                     := '0';

    ------ Register signals (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit
    signal regs_read_arr        : t_std32_array(IPB_TTC_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(IPB_TTC_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(IPB_TTC_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(IPB_TTC_NUM_REGS - 1 downto 0);
    signal regs_read_pulse_arr  : std_logic_vector(IPB_TTC_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(IPB_TTC_NUM_REGS - 1 downto 0);
    ------ End of register signals
    
--============================================================================
--                                                          Architecture begin
--============================================================================

begin
    i_reset_sync: 
    entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => clk_40,
            sync_o  => reset
        );

    i_ttc_clocks:
    entity work.ttc_clocks
        port map(
            clk_40_ttc_p_i       => clk_40_ttc_p_i,
            clk_40_ttc_n_i       => clk_40_ttc_n_i,
            mmcm_rst_i           => ttc_ctrl.mmcm_reset,
            mmcm_locked_o        => ttc_stat.mmcm_locked,
            ttc_mmcm_ps_clk_i    => clk_40,
            ttc_mmcm_ps_clk_en_i => ttc_ctrl.mmcm_phase_shift,
            clk_40_bufg_o        => clk_40,
            clk_80_bufg_o        => clk_80,
            clk_160_bufg_o       => clk_160,
            clk_240_bufg_o       => clk_240,
            clk_320_bufg_o       => clk_320
        );

    i_ttc_cmd:
    entity work.ttc_cmd
        port map(
            clk_40_i             => clk_40,
            ttc_data_p_i         => ttc_data_p_i,
            ttc_data_n_i         => ttc_data_n_i,
            ttc_cmd_o            => ttc_cmd,
            ttc_l1a_o            => ttc_l1a,
            tcc_err_cnt_rst_i    => ttc_ctrl_i.stat_reset or reset,
            ttc_err_single_cnt_o => ttc_status.single_err,
            ttc_err_double_cnt_o => ttc_status.double_err
        );

    p_cmd:
    process(clk_40) is
    begin
        if (rising_edge(clk_40)) then
            if (reset = '1') then
                bc0_cmd        <= '0';
                ec0_cmd        <= '0';
                resync_cmd     <= '0';
                oc0_cmd        <= '0';
                start_cmd      <= '0';
                stop_cmd       <= '0';
                test_sync_cmd  <= '0';
                hard_reset_cmd <= '0';
                calpulse_cmd   <= '0';
                l1a_cmd        <= '0';
            else
                if (ttc_cmd = ttc_conf.cmd_bc0) then
                    bc0_cmd <= '1';
                else
                    bc0_cmd <= '0';
                end if;
                if (ttc_cmd = ttc_conf.cmd_ec0) then
                    ec0_cmd <= '1';
                else
                    ec0_cmd <= '0';
                end if;
                if (ttc_cmd = ttc_conf.cmd_resync) then
                    resync_cmd <= '1';
                else
                    resync_cmd <= '0';
                end if;
                if (ttc_cmd = ttc_conf.cmd_oc0) then
                    oc0_cmd <= '1';
                else
                    oc0_cmd <= '0';
                end if;
                if (ttc_cmd = ttc_conf.cmd_hard_reset) then
                    s_hart_reset_cmd <= '1';
                else
                    hard_reset_cmd <= '0';
                end if;
                if (ttc_cmd = ttc_conf.cmd_calpulse) then
                    calpulse_cmd <= '1';
                else
                    calpulse_cmd <= '0';
                end if;
                if (ttc_cmd = ttc_conf.cmd_start) then
                    start_cmd <= '1';
                else
                    start_cmd <= '0';
                end if;
                if (ttc_cmd = ttc_conf.cmd_stop) then
                    stop_cmd <= '1';
                else
                    stop_cmd <= '0';
                end if;
                if (ttc_cmd = ttc_conf.cmd_test_sync) then
                    test_sync_cmd <= '1';
                else
                    test_sync_cmd <= '0';
                end if;

                l1a_cmd <= ttc_l1a and ttc_ctrl.l1a_enable;

            end if;

        end if;
    end process p_cmd;

    p_orbit_cnt:
    process(clk_40) is
    begin
        if (rising_edge(clk_40)) then
            if (reset = '1') then
                orbit_cnt <= (others => '0');
            else
                if (oc0_cmd = '1') then
                    orbit_cnt <= (others => '0');
                elsif (bc0_cmd = '1') then
                    orbit_cnt <= std_logic_vector(unsigned(orbit_cnt) + 1);
                end if;
            end if;

        end if;
    end process p_orbit_cnt;

    p_l1id_cnt:
    process(clk_40) is
    begin
        if (rising_edge(clk_40)) then
            if (reset = '1') then
                l1id_cnt <= (others => '0');
            else
                if (ec0_cmd = '1') then
                    l1id_cnt <= (others => '0');
                elsif (l1a_cmd = '1') then
                    l1id_cnt <= std_logic_vector(unsigned(l1id_cnt) + 1);
                end if;
            end if;

        end if;
    end process p_l1id_cnt;

    p_bx_cnt:
    process(clk_40) is
    begin
        if (rising_edge(clk_40)) then
            if (reset = '1') then
                bc0_cmd <= (others => '0');
            else
                if (bc0_cmd = '1') then
                    s_bc_cnt <= (others => '0');
                else
                    bx_cnt <= std_logic_vector(unsigned(bx_cnt) + 1);
                end if;
            end if;

        end if;
    end process bx_cnt;

    p_mini_spy:
    process(clk_40) is
    begin
        if rising_edge(clk) then
            if rst = '1' then
            else
            end if;
        end if;
    end process mini_spy;

    ttc_daq_cntrs_o.orbit <= orbit_cnt;
    ttc_daq_cntrs_o.l1id  <= l1id_cnt;
    ttc_daq_cntrs_o.bx    <= bx_cnt;

    ttc_cmds_arr(0) <= l1a_cmd;
    ttc_cmds_arr(1) <= bc0_cmd;
    ttc_cmds_arr(2) <= ec0_cmd;
    ttc_cmds_arr(3) <= resync_cmd;
    ttc_cmds_arr(4) <= oc0_cmd;
    ttc_cmds_arr(5) <= hard_reset_cmd;
    ttc_cmds_arr(6) <= calpulse_cmd;
    ttc_cmds_arr(7) <= start_cmd;
    ttc_cmds_arr(8) <= stop_cmd;
    ttc_cmds_arr(9) <= test_sync_cmd;

    gen_ttc_cmd_cnt:
    for i in 0 to C_NUM_OF_DECODED_TTC_CMDS - 1 generate
        process(clk_40) is
        begin
            if (rising_edge(clk_40)) then
                if (ttc_ctrl.stat_reset = '1' or reset = '1') then
                    ttc_cmds_cnt_arr(i) <= (others => '0');
                elsif (ttc_cmds_arr(i) = '1') then
                    ttc_cmds_cnt_arr(i) <= std_logic_vector(unsigned(ttc_cmds_cnt_arr(i)) + 1);
                end if;
            end if;
        end process;
    end generate;

    ttc_cmds_o.l1a        <= l1a_cmd;
    ttc_cmds_o.bc0        <= bc0_cmd;
    ttc_cmds_o.ec0        <= ec0_cmd;
    ttc_cmds_o.resync     <= resync_cmd;
    ttc_cmds_o.hard_reset <= hard_reset_cmd;
    ttc_cmds_o.calpulse   <= calpulse_cmd;
    ttc_cmds_o.start      <= start_cmd;
    ttc_cmds_o.stop       <= stop_cmd;
    ttc_cmds_o.test_sync  <= test_sync_cmd;

    ttc_clks_o.clk_40  <= clk_40;
    ttc_clks_o.clk_80  <= clk_80;
    ttc_clks_o.clk_160 <= clk_160;
    ttc_clks_o.clk_240 <= clk_240;
    ttc_clks_o.clk_320 <= clk_320;

    --==== Registers ================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --===============================================================================================
    
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
            g_NUM_REGS             => IPB_TTC_NUM_REGS,
            g_ADDR_HIGH_BIT        => g_ADDR_HIGH_BIT,
            g_ADDR_LOW_BIT         => g_ADDR_LOW_BIT,
            g_USE_INDIVIDUAL_ADDRS => "FALSE"
        )
        port map(
            ipb_reset_i            => ipb_reset_i,
            ipb_clk_i              => ipb_clk_i,
            ipb_mosi_i             => ipb_mosi_i,
            ipb_miso_o             => ipb_miso_o,
            usr_clk_i              => clk_40,
            regs_read_arr_i        => regs_read_arr,
            regs_write_arr_o       => regs_write_arr,
            read_pulse_arr_o       => regs_read_pulse_arr,
            write_pulse_arr_o      => regs_write_pulse_arr,
            individual_addrs_arr_i => regs_addresses,
            regs_defaults_arr_i    => regs_defaults
        );

    --==== End of registers =========================================================================

end ttc_arch;
--============================================================================
--                                                            Architecture end
--============================================================================

-------------------------------------------------------------------------------
--                                                                            
--       Unit Name: gth_wrapper                                            
--                                                                            
--     Description: 
--
--                                                                            
-------------------------------------------------------------------------------
--                                                                            
--           Notes:                                                           
--                                                                            
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use ieee.std_logic_misc.all;

library UNISIM;
use UNISIM.VCOMPONENTS.all;

library work;
use work.gth_pkg.all;
use work.gem_pkg.all;

use work.system_package.all;

--============================================================================
--                                                          Entity declaration
--============================================================================
entity gth_wrapper is
  generic
    (
      g_EXAMPLE_SIMULATION     : integer                := 0;
      g_STABLE_CLOCK_PERIOD    : integer range 4 to 250 := 20;  --Period of the stable clock driving this state-machine, unit is [ns]
      g_NUM_OF_GTH_GTs         : integer                := 64;
      g_NUM_OF_GTH_COMMONs     : integer                := 16;
      g_GT_SIM_GTRESET_SPEEDUP : string                 := "FALSE"  -- Set to "TRUE" to speed up sim reset

      );
  port (

    clk_stable_i : in std_logic;

    refclk_F_0_p_i : in std_logic_vector (3 downto 0);
    refclk_F_0_n_i : in std_logic_vector (3 downto 0);
    refclk_F_1_p_i : in std_logic_vector (3 downto 0);
    refclk_F_1_n_i : in std_logic_vector (3 downto 0);
    refclk_B_0_p_i : in std_logic_vector (3 downto 1);
    refclk_B_0_n_i : in std_logic_vector (3 downto 1);
    refclk_B_1_p_i : in std_logic_vector (3 downto 1);
    refclk_B_1_n_i : in std_logic_vector (3 downto 1);

    clk_gth_tx_usrclk_arr_o : out std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
    clk_gth_rx_usrclk_arr_o : out std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);

    ------------------------

    gth_cpll_status_arr_o : out t_gth_cpll_status_arr(g_NUM_OF_GTH_GTs-1 downto 0);

    ------------------------
    -- GTH common

    gth_common_reset_i      : in  std_logic_vector(g_NUM_OF_GTH_COMMONs-1 downto 0);
    gth_common_status_arr_o : out t_gth_common_status_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);

    gth_common_drp_arr_i : in  t_gth_common_drp_in_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);
    gth_common_drp_arr_o : out t_gth_common_drp_out_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);
    ------------------------

    gth_gt_txreset_i : in std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
    gth_gt_rxreset_i : in std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);

    gth_gt_txreset_done_o : out std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
    gth_gt_rxreset_done_o : out std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);

    gth_rx_serial_arr_i : in  t_gth_rx_serial_arr(g_NUM_OF_GTH_GTs-1 downto 0);
    gth_tx_serial_arr_o : out t_gth_tx_serial_arr(g_NUM_OF_GTH_GTs-1 downto 0);

    gth_gt_drp_arr_i : in  t_gth_gt_drp_in_arr(g_NUM_OF_GTH_GTs-1 downto 0);
    gth_gt_drp_arr_o : out t_gth_gt_drp_out_arr(g_NUM_OF_GTH_GTs-1 downto 0);

    gth_tx_ctrl_arr_i   : in  t_gth_tx_ctrl_arr(g_NUM_OF_GTH_GTs-1 downto 0);
    gth_tx_status_arr_o : out t_gth_tx_status_arr(g_NUM_OF_GTH_GTs-1 downto 0);

    gth_rx_ctrl_arr_i   : in t_gth_rx_ctrl_arr(g_NUM_OF_GTH_GTs-1 downto 0);
    gth_rx_ctrl_2_arr_i : in t_gth_rx_ctrl_2_arr(g_NUM_OF_GTH_GTs-1 downto 0);

    gth_rx_status_arr_o : out t_gth_rx_status_arr(g_NUM_OF_GTH_GTs-1 downto 0);

    gth_misc_ctrl_arr_i   : in  t_gth_misc_ctrl_arr(g_NUM_OF_GTH_GTs-1 downto 0);
    gth_misc_status_arr_o : out t_gth_misc_status_arr(g_NUM_OF_GTH_GTs-1 downto 0);

    gth_tx_data_arr_i : in  t_gt_8b10b_tx_data_arr(g_NUM_OF_GTH_GTs-1 downto 0);
    gth_rx_data_arr_o : out t_gt_8b10b_rx_data_arr(g_NUM_OF_GTH_GTs-1 downto 0)
    );
end gth_wrapper;

--============================================================================
--                                                        Architecture section
--============================================================================
architecture gth_wrapper_arch of gth_wrapper is

--============================================================================
--                                                         Signal declarations
--============================================================================

  signal s_refclk_F_0 : std_logic_vector (3 downto 0);
  signal s_refclk_F_1 : std_logic_vector (3 downto 0);
  signal s_refclk_B_0 : std_logic_vector (3 downto 1);
  signal s_refclk_B_1 : std_logic_vector (3 downto 1);

  attribute syn_noclockbuf : boolean;

  attribute syn_noclockbuf of s_refclk_F_0 : signal is true;
  attribute syn_noclockbuf of s_refclk_F_1 : signal is true;
  attribute syn_noclockbuf of s_refclk_B_0 : signal is true;
  attribute syn_noclockbuf of s_refclk_B_1 : signal is true;


  signal s_gth_rx_serial_arr : t_gth_rx_serial_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_tx_serial_arr : t_gth_tx_serial_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_gt_clk_in_arr  : t_gth_gt_clk_in_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_gt_clk_out_arr : t_gth_gt_clk_out_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_cpll_ctrl_arr   : t_gth_cpll_ctrl_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_cpll_init_arr   : t_gth_cpll_init_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_cpll_status_arr : t_gth_cpll_status_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_gt_drp_in_arr  : t_gth_gt_drp_in_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_gt_drp_out_arr : t_gth_gt_drp_out_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_tx_ctrl_arr   : t_gth_tx_ctrl_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_tx_init_arr   : t_gth_tx_init_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_tx_status_arr : t_gth_tx_status_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_rx_ctrl_arr   : t_gth_rx_ctrl_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_rx_ctrl_2_arr : t_gth_rx_ctrl_2_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_rx_init_arr : t_gth_rx_init_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_rx_status_arr : t_gth_rx_status_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_misc_ctrl_arr   : t_gth_misc_ctrl_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_misc_status_arr : t_gth_misc_status_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_tx_data_arr : t_gt_8b10b_tx_data_arr(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_rx_data_arr : t_gt_8b10b_rx_data_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  ---------------------

  signal s_gth_common_clk_in_arr  : t_gth_common_clk_in_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);
  signal s_gth_common_clk_out_arr : t_gth_common_clk_out_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);

  signal s_gth_common_ctrl_arr   : t_gth_common_ctrl_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);
  signal s_gth_common_status_arr : t_gth_common_status_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);

  signal s_gth_common_drp_in_arr  : t_gth_common_drp_in_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);
  signal s_gth_common_drp_out_arr : t_gth_common_drp_out_arr(g_NUM_OF_GTH_COMMONs-1 downto 0);

  ---------------------
  function get_cdrlock_time(is_sim : in integer) return integer is
    variable lock_time : integer;
  begin
    if (is_sim = 1) then
      lock_time := 1000;
    else
      lock_time := 50000 / integer(3.2);  --Typical CDR lock time is 50,000UI as per DS183
    end if;
    return lock_time;
  end function;

  constant C_RX_CDRLOCK_TIME   : integer := get_cdrlock_time(g_EXAMPLE_SIMULATION);  -- 200us
  constant C_WAIT_TIME_CDRLOCK : integer := C_RX_CDRLOCK_TIME / g_STABLE_CLOCK_PERIOD;  -- 200 us time-out

  type t_rx_cdr_lock_counter_arr is array(integer range <>) of integer range 0 to C_WAIT_TIME_CDRLOCK;

  signal s_gth_tx_run_phalignment      : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_tx_run_phalignment_done : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_tx_rst_phalignment      : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_rx_run_phalignment      : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_rx_run_phalignment_done : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_rx_rst_phalignment      : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_gth_recclk_stable      : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_rx_cdrlocked       : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_gth_rx_cdrlock_counter : t_rx_cdr_lock_counter_arr(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_clk_gth_tx_usrclk_arr : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_clk_gth_rx_usrclk_arr : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);

  signal s_tx_startup_fsm_mmcm_reset : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0);
  signal s_tx_startup_fsm_mmcm_lock  : std_logic_vector(g_NUM_OF_GTH_GTs-1 downto 0) := (others => '1');


  signal s_GTH_4p8g_TX_MMCM_reset  : std_logic;
  signal s_GTH_4p8g_TX_MMCM_locked : std_logic;


--============================================================================
--                                                          Architecture begin
--============================================================================

begin

  gen_tx_mmcm_sigs : for n in 0 to g_NUM_OF_GTH_GTs-1 generate


    gen_gth_4p8g_txuserclk : if c_gth_config_arr(n).gth_link_type = gth_4p8g generate

      gen_gth_4p8g_txuserclk_master : if c_gth_config_arr(n).gth_txclk_out_master = true generate

        s_GTH_4p8g_TX_MMCM_reset <= s_tx_startup_fsm_mmcm_reset(n);

        s_tx_startup_fsm_mmcm_lock(n) <= s_GTH_4p8g_TX_MMCM_locked;

      end generate;
    end generate;
  end generate;

  i_gth_clk_bufs : entity work.gth_clk_bufs
    generic map
    (
      g_NUM_OF_GTH_GTs => g_NUM_OF_GTH_GTs
      )
    port map
    (

      GTH_4p8g_TX_MMCM_reset_i  => s_GTH_4p8g_TX_MMCM_reset,
      GTH_4p8g_TX_MMCM_locked_o => s_GTH_4p8g_TX_MMCM_locked,

      refclk_F_0_p_i => refclk_F_0_p_i,
      refclk_F_0_n_i => refclk_F_0_n_i,
      refclk_F_1_p_i => refclk_F_1_p_i,
      refclk_F_1_n_i => refclk_F_1_n_i,
      refclk_B_0_p_i => refclk_B_0_p_i,
      refclk_B_0_n_i => refclk_B_0_n_i,
      refclk_B_1_p_i => refclk_B_1_p_i,
      refclk_B_1_n_i => refclk_B_1_n_i,

      refclk_F_0_o => s_refclk_F_0,
      refclk_F_1_o => s_refclk_F_1,
      refclk_B_0_o => s_refclk_B_0,
      refclk_B_1_o => s_refclk_B_1,

      gth_gt_clk_out_arr_i => s_gth_gt_clk_out_arr,

      clk_gth_tx_usrclk_arr_o => s_clk_gth_tx_usrclk_arr,
      clk_gth_rx_usrclk_arr_o => s_clk_gth_rx_usrclk_arr

      );

  clk_gth_tx_usrclk_arr_o <= s_clk_gth_tx_usrclk_arr;
  clk_gth_rx_usrclk_arr_o <= s_clk_gth_rx_usrclk_arr;

------------------------

  gen_qpll_refclk_assign_Q110_to_Q111 : for i in 0 to 1 generate
  begin
    gen_qpll_inner : for j in 0 to 3 generate
    begin
      s_gth_gt_clk_in_arr(i*4+j).GTREFCLK0  <= s_refclk_F_0(3);
      s_gth_gt_clk_in_arr(i*4+j).qpllclk    <= s_gth_common_clk_out_arr(i).QPLLCLK;
      s_gth_gt_clk_in_arr(i*4+j).qpllrefclk <= s_gth_common_clk_out_arr(i).QPLLREFCLK;
    end generate;
  end generate;

  gen_qpll_refclk_assign_Q112_to_Q114 : for i in 2 to 4 generate
  begin
    gen_qpll_inner : for j in 0 to 3 generate
    begin
      s_gth_gt_clk_in_arr(i*4+j).GTREFCLK0  <= s_refclk_F_0(2);
      s_gth_gt_clk_in_arr(i*4+j).qpllclk    <= s_gth_common_clk_out_arr(i).QPLLCLK;
      s_gth_gt_clk_in_arr(i*4+j).qpllrefclk <= s_gth_common_clk_out_arr(i).QPLLREFCLK;
    end generate;
  end generate;

  gen_qpll_refclk_assign_Q115_to_Q117 : for i in 5 to 7 generate
  begin
    gen_qpll_inner : for j in 0 to 3 generate
    begin
      s_gth_gt_clk_in_arr(i*4+j).GTREFCLK0  <= s_refclk_F_0(1);
      s_gth_gt_clk_in_arr(i*4+j).qpllclk    <= s_gth_common_clk_out_arr(i).QPLLCLK;
      s_gth_gt_clk_in_arr(i*4+j).qpllrefclk <= s_gth_common_clk_out_arr(i).QPLLREFCLK;
    end generate;
  end generate;

  gen_qpll_refclk_assign_Q118 : for i in 8 to 8 generate
  begin
    gen_qpll_inner : for j in 0 to 3 generate
    begin
      s_gth_gt_clk_in_arr(i*4+j).GTREFCLK0  <= s_refclk_F_0(0);
      s_gth_gt_clk_in_arr(i*4+j).qpllclk    <= s_gth_common_clk_out_arr(i).QPLLCLK;
      s_gth_gt_clk_in_arr(i*4+j).qpllrefclk <= s_gth_common_clk_out_arr(i).QPLLREFCLK;
    end generate;
  end generate;

--------

  s_gth_rx_serial_arr <= gth_rx_serial_arr_i;
  gth_tx_serial_arr_o <= s_gth_tx_serial_arr;

  s_gth_gt_drp_in_arr <= gth_gt_drp_arr_i;
  gth_gt_drp_arr_o    <= s_gth_gt_drp_out_arr;

  s_gth_tx_ctrl_arr     <= gth_tx_ctrl_arr_i;
  gth_tx_status_arr_o   <= s_gth_tx_status_arr;
  s_gth_rx_ctrl_arr     <= gth_rx_ctrl_arr_i;
  s_gth_rx_ctrl_2_arr   <= gth_rx_ctrl_2_arr_i;
  gth_rx_status_arr_o   <= s_gth_rx_status_arr;
  s_gth_misc_ctrl_arr   <= gth_misc_ctrl_arr_i;
  gth_misc_status_arr_o <= s_gth_misc_status_arr;


  gen_gth_single : for n in 0 to (g_NUM_OF_GTH_GTs-1) generate
  begin

-- From Xilinx UG476
-- The CPLLREFCLKSEL port is required when multiple reference clock sources are 
-- connected to this multiplexer. A single reference clock is most commonly used. 
-- In this case, the CPLLREFCLKSEL port can be tied to 3'b001, and the Xilinx software 
-- tools handle the complexity of the multiplexers and associated routing.
    s_gth_cpll_ctrl_arr(n).CPLLREFCLKSEL  <= "001";  -- Let the tool figure out proper reference clock routing
    s_gth_cpll_ctrl_arr(n).cplllockdetclk <= clk_stable_i;

    s_gth_gt_clk_in_arr(n).rxusrclk  <= s_clk_gth_rx_usrclk_arr(n);
    s_gth_gt_clk_in_arr(n).rxusrclk2 <= s_clk_gth_rx_usrclk_arr(n);
    s_gth_gt_clk_in_arr(n).txusrclk  <= s_clk_gth_tx_usrclk_arr(n);
    s_gth_gt_clk_in_arr(n).txusrclk2 <= s_clk_gth_tx_usrclk_arr(n);


    gen_gth_3p2g : if c_gth_config_arr(n).gth_link_type = gth_3p2g generate

      s_gth_tx_data_arr(n) <= gth_tx_data_arr_i(n);
      gth_rx_data_arr_o(n) <= s_gth_rx_data_arr(n);
      s_gth_rx_status_arr(n).rxnotintable <= s_gth_rx_data_arr(n).rxnotintable;
      s_gth_rx_status_arr(n).rxdisperr <= s_gth_rx_data_arr(n).rxdisperr;

      i_gth_single_3p2g : entity work.gth_single_3p2g
        generic map
        (
                                        -- Simulation attributes
          g_GT_SIM_GTRESET_SPEEDUP => g_GT_SIM_GTRESET_SPEEDUP
          )
        port map
        (
          gth_rx_serial_i => s_gth_rx_serial_arr(n),
          gth_tx_serial_o => s_gth_tx_serial_arr(n),
          gth_gt_clk_i    => s_gth_gt_clk_in_arr(n),
          gth_gt_clk_o    => s_gth_gt_clk_out_arr(n),

          gth_cpll_ctrl_i   => s_gth_cpll_ctrl_arr(n),
          gth_cpll_init_i   => s_gth_cpll_init_arr(n),
          gth_cpll_status_o => s_gth_cpll_status_arr(n),

          gth_gt_drp_i      => s_gth_gt_drp_in_arr(n),
          gth_gt_drp_o      => s_gth_gt_drp_out_arr(n),
          gth_tx_ctrl_i     => s_gth_tx_ctrl_arr(n),
          gth_tx_init_i     => s_gth_tx_init_arr(n),
          gth_tx_status_o   => s_gth_tx_status_arr(n),
          gth_rx_ctrl_i     => s_gth_rx_ctrl_arr(n),
          gth_rx_ctrl_2_i   => s_gth_rx_ctrl_2_arr(n),
          gth_rx_init_i     => s_gth_rx_init_arr(n),
          gth_rx_status_o   => s_gth_rx_status_arr(n),
          gth_misc_ctrl_i   => s_gth_misc_ctrl_arr(n),
          gth_misc_status_o => s_gth_misc_status_arr(n),
          gth_tx_data_i     => s_gth_tx_data_arr(n),
          gth_rx_data_o     => s_gth_rx_data_arr(n)
          );
        
    end generate;


    gen_gth_4p8g : if c_gth_config_arr(n).gth_link_type = gth_4p8g generate

      -------------  GT txdata_i Assignments for 20 bit datapath  -------  
      s_gth_tx_data_arr(n).txdata <= x"0000" &
                                     gth_tx_data_arr_i(n).txdata(17 downto 10) &
                                     gth_tx_data_arr_i(n).txdata(7 downto 0);

      s_gth_tx_data_arr(n).txchardispmode <= "00" &
                                             gth_tx_data_arr_i(n).txdata(19) &
                                             gth_tx_data_arr_i(n).txdata(9);

      s_gth_tx_data_arr(n).txchardispval <= "00" &
                                            gth_tx_data_arr_i(n).txdata(18) &
                                            gth_tx_data_arr_i(n).txdata(8);

      s_gth_tx_data_arr(n).txcharisk <= gth_tx_data_arr_i(n).txcharisk;

      -------------  GT RXDATA Assignments for 20 bit datapath  -------  

      gth_rx_data_arr_o(n).rxdata <= x"000" &
                                     s_gth_rx_data_arr(n).rxdisperr(1) &
                                     s_gth_rx_data_arr(n).rxcharisk(1) &
                                     s_gth_rx_data_arr(n).rxdata(15 downto 8) &
                                     s_gth_rx_data_arr(n).rxdisperr(0) &
                                     s_gth_rx_data_arr(n).rxcharisk(0) &
                                     s_gth_rx_data_arr(n).rxdata(7 downto 0);


      gth_rx_data_arr_o(n).rxbyteisaligned <= s_gth_rx_data_arr(n).rxbyteisaligned;
      gth_rx_data_arr_o(n).rxbyterealign   <= s_gth_rx_data_arr(n).rxbyterealign;
      gth_rx_data_arr_o(n).rxcommadet      <= s_gth_rx_data_arr(n).rxcommadet;
      gth_rx_data_arr_o(n).rxdisperr       <= s_gth_rx_data_arr(n).rxdisperr;
      gth_rx_data_arr_o(n).rxnotintable    <= s_gth_rx_data_arr(n).rxnotintable;
      gth_rx_data_arr_o(n).rxchariscomma   <= s_gth_rx_data_arr(n).rxchariscomma;
      gth_rx_data_arr_o(n).rxcharisk       <= s_gth_rx_data_arr(n).rxcharisk;

      i_gth_single_4p8g : entity work.gth_single_4p8g
        generic map
        (
                                        -- Simulation attributes
          g_GT_SIM_GTRESET_SPEEDUP => g_GT_SIM_GTRESET_SPEEDUP
          )
        port map
        (
          gth_rx_serial_i => s_gth_rx_serial_arr(n),
          gth_tx_serial_o => s_gth_tx_serial_arr(n),
          gth_gt_clk_i    => s_gth_gt_clk_in_arr(n),
          gth_gt_clk_o    => s_gth_gt_clk_out_arr(n),

          gth_cpll_ctrl_i   => s_gth_cpll_ctrl_arr(n),
          gth_cpll_init_i   => s_gth_cpll_init_arr(n),
          gth_cpll_status_o => s_gth_cpll_status_arr(n),

          gth_gt_drp_i      => s_gth_gt_drp_in_arr(n),
          gth_gt_drp_o      => s_gth_gt_drp_out_arr(n),
          gth_tx_ctrl_i     => s_gth_tx_ctrl_arr(n),
          gth_tx_init_i     => s_gth_tx_init_arr(n),
          gth_tx_status_o   => s_gth_tx_status_arr(n),
          gth_rx_ctrl_i     => s_gth_rx_ctrl_arr(n),
          gth_rx_ctrl_2_i   => s_gth_rx_ctrl_2_arr(n),
          gth_rx_init_i     => s_gth_rx_init_arr(n),
          gth_rx_status_o   => s_gth_rx_status_arr(n),
          gth_misc_ctrl_i   => s_gth_misc_ctrl_arr(n),
          gth_misc_status_o => s_gth_misc_status_arr(n),
          gth_tx_data_i     => s_gth_tx_data_arr(n),
          gth_rx_data_o     => s_gth_rx_data_arr(n)
          );

    end generate;
  end generate;


  s_gth_common_drp_in_arr <= gth_common_drp_arr_i;
  gth_common_drp_arr_o    <= s_gth_common_drp_out_arr;

  s_gth_common_clk_in_arr(0).GTREFCLK0 <= s_refclk_F_1(3);
  s_gth_common_clk_in_arr(1).GTREFCLK0 <= s_refclk_F_1(3);

  s_gth_common_clk_in_arr(2).GTREFCLK0 <= s_refclk_F_1(2);
  s_gth_common_clk_in_arr(3).GTREFCLK0 <= s_refclk_F_1(2);
  s_gth_common_clk_in_arr(4).GTREFCLK0 <= s_refclk_F_1(2);

  s_gth_common_clk_in_arr(5).GTREFCLK0 <= s_refclk_F_1(1);
  s_gth_common_clk_in_arr(6).GTREFCLK0 <= s_refclk_F_1(1);
  s_gth_common_clk_in_arr(7).GTREFCLK0 <= s_refclk_F_1(1);

  s_gth_common_clk_in_arr(8).GTREFCLK0 <= s_refclk_F_1(0);
  s_gth_common_clk_in_arr(9).GTREFCLK0 <= s_refclk_F_1(0);


  s_gth_common_clk_in_arr(10).GTREFCLK0 <= s_refclk_B_1(3);
  s_gth_common_clk_in_arr(11).GTREFCLK0 <= s_refclk_B_1(3);

  s_gth_common_clk_in_arr(12).GTREFCLK0 <= s_refclk_B_1(2);
  s_gth_common_clk_in_arr(13).GTREFCLK0 <= s_refclk_B_1(2);
  s_gth_common_clk_in_arr(14).GTREFCLK0 <= s_refclk_B_1(2);

  s_gth_common_clk_in_arr(15).GTREFCLK0 <= s_refclk_B_1(1);

  gth_common_status_arr_o <= s_gth_common_status_arr;
  gth_cpll_status_arr_o   <= s_gth_cpll_status_arr;


  -- GTH Common not used in this demo project for TAMU. Commented out.
  gen_gth_common : for n in 0 to (g_NUM_OF_GTH_COMMONs-1) generate
  begin

    s_gth_common_ctrl_arr(n).QPLLRESET <= gth_common_reset_i(n);

    -- From Xilinx UG476
    -- The QPLLREFCLKSEL port is required when multiple reference clock sources are 
    -- connected to this multiplexer. A single reference clock is most commonly used. 
    -- In this case, the QPLLREFCLKSEL port can be tied to 3'b001, and the Xilinx software 
    -- tools handle the complexity of the multiplexers and associated routing.
    s_gth_common_ctrl_arr(n).QPLLREFCLKSEL <= "001";  -- Let the tool figure out proper reference clock routing

--    i_gth_common : entity work.gth_common
--      generic map
--      (
--                                        -- Simulation attributes
--        g_GT_SIM_GTRESET_SPEEDUP => g_GT_SIM_GTRESET_SPEEDUP,  -- Set to "true" to speed up sim reset
--        g_STABLE_CLOCK_PERIOD    => g_STABLE_CLOCK_PERIOD  -- Period of the stable clock driving this state-machine, unit is [ns]
--        )
--      port map
--      (
--        clk_stable_i        => clk_stable_i,
--        gth_common_clk_i    => s_gth_common_clk_in_arr(n),
--        gth_common_clk_o    => s_gth_common_clk_out_arr(n),
--        gth_common_ctrl_i   => s_gth_common_ctrl_arr(n),
--        gth_common_status_o => s_gth_common_status_arr(n),
--        gth_common_drp_i    => s_gth_common_drp_in_arr(n),
--        gth_common_drp_o    => s_gth_common_drp_out_arr(n)
--        );

  end generate;

  gen_gt_resetfsm : for i in 0 to (g_NUM_OF_GTH_GTs/4-1) generate
  begin
    gen_txresetfsm_inner : for j in 0 to 3 generate
    begin

      i_gt_txresetfsm : entity work.gth_single_TX_STARTUP_FSM

        generic map(
          EXAMPLE_SIMULATION     => g_EXAMPLE_SIMULATION,
          STABLE_CLOCK_PERIOD    => g_STABLE_CLOCK_PERIOD,  -- Period of the stable clock driving this state-machine, unit is [ns]
          RETRY_COUNTER_BITWIDTH => 8,
          TX_QPLL_USED           => false,  -- the TX and RX Reset FSMs must
          RX_QPLL_USED           => false,  -- share these two generic values
          PHASE_ALIGNMENT_MANUAL => true  -- Decision if a manual phase-alignment is necessary or the automatic
                                          -- is enough. For single-lane applications the automatic alignment is
                                          -- sufficient
          )
        port map (
          STABLE_CLOCK      => clk_stable_i,
          TXUSERCLK         => s_clk_gth_tx_usrclk_arr(i*4+j),
          SOFT_RESET        => gth_gt_txreset_i(i*4+j),
          QPLLREFCLKLOST    => '0',
          CPLLREFCLKLOST    => '0',
          QPLLLOCK          => '1',
          CPLLLOCK          => s_gth_cpll_status_arr(i).CPLLLOCK,
          TXRESETDONE       => s_gth_tx_status_arr(i*4+j).txresetdone,
          MMCM_LOCK         => s_tx_startup_fsm_mmcm_lock(i*4+j),
          GTTXRESET         => s_gth_tx_init_arr(i*4+j).gttxreset,
          MMCM_RESET        => s_tx_startup_fsm_mmcm_reset(i*4+j),
          QPLL_RESET        => open,
          CPLL_RESET        => open,
          TX_FSM_RESET_DONE => gth_gt_txreset_done_o(i*4+j),
          TXUSERRDY         => s_gth_tx_init_arr(i*4+j).txuserrdy,
          RUN_PHALIGNMENT   => s_gth_tx_run_phalignment(i*4+j),
          RESET_PHALIGNMENT => s_gth_tx_rst_phalignment(i*4+j),
          PHALIGNMENT_DONE  => s_gth_tx_run_phalignment_done(i*4+j),
          RETRY_COUNTER     => open
          );

      i_gt_rxresetfsm : entity work.gth_single_RX_STARTUP_FSM

        generic map(
          EXAMPLE_SIMULATION     => g_EXAMPLE_SIMULATION,
          EQ_MODE                => "LPM",  --Rx Equalization Mode - Set to DFE or LPM
          STABLE_CLOCK_PERIOD    => g_STABLE_CLOCK_PERIOD,  --Period of the stable clock driving this state-machine, unit is [ns]
          RETRY_COUNTER_BITWIDTH => 8,
          TX_QPLL_USED           => false,  -- the TX and RX Reset FSMs must
          RX_QPLL_USED           => false,  -- share these two generic values
          PHASE_ALIGNMENT_MANUAL => false  -- Decision if a manual phase-alignment is necessary or the automatic
                                           -- is enough. For single-lane applications the automatic alignment is
                                           -- sufficient
          )
        port map (
          STABLE_CLOCK             => clk_stable_i,
          RXUSERCLK                => s_clk_gth_rx_usrclk_arr(i*4+j),
          SOFT_RESET               => gth_gt_rxreset_i(i*4+j),
          DONT_RESET_ON_DATA_ERROR => '1',
          RXPMARESETDONE           => s_gth_rx_status_arr(i*4+j).RXPMARESETDONE,
          RXOUTCLK                 => s_gth_gt_clk_out_arr(i*4+j).rxoutclk,
          QPLLREFCLKLOST           => '0',
          CPLLREFCLKLOST           => s_gth_cpll_status_arr(i).CPLLREFCLKLOST,
          QPLLLOCK                 => '1',
          CPLLLOCK                 => s_gth_cpll_status_arr(i).CPLLLOCK,
          RXRESETDONE              => s_gth_rx_status_arr(i*4+j).rxresetdone,
          MMCM_LOCK                => '1',
          RECCLK_STABLE            => s_gth_recclk_stable(i*4+j),
          RECCLK_MONITOR_RESTART   => '0',
          DATA_VALID               => '1',
          TXUSERRDY                => '1',
          GTRXRESET                => s_gth_rx_init_arr(i*4+j).gtrxreset,
          MMCM_RESET               => open,
          QPLL_RESET               => open,
          CPLL_RESET               => s_gth_cpll_init_arr(i*4+j).cpllreset,
          RX_FSM_RESET_DONE        => gth_gt_rxreset_done_o(i*4+j),
          RXUSERRDY                => s_gth_rx_init_arr(i*4+j).rxuserrdy,
          RUN_PHALIGNMENT          => s_gth_rx_run_phalignment(i*4+j),
          RESET_PHALIGNMENT        => s_gth_rx_rst_phalignment(i*4+j),
          PHALIGNMENT_DONE         => s_gth_rx_run_phalignment_done(i*4+j),
          RXDFEAGCHOLD             => s_gth_rx_init_arr(i*4+j).RXDFEAGCHOLD,
          RXDFELFHOLD              => s_gth_rx_init_arr(i*4+j).RXDFELFHOLD,
          RXLPMLFHOLD              => s_gth_rx_init_arr(i*4+j).RXLPMLFHOLD,
          RXLPMHFHOLD              => s_gth_rx_init_arr(i*4+j).RXLPMHFHOLD,
          RETRY_COUNTER            => open
          );

      s_gth_rx_init_arr(i*4+j).rxdfeagcovrden  <= '0';
      s_gth_rx_init_arr(i*4+j).rxdfelpmreset   <= '0';
      s_gth_rx_init_arr(i*4+j).rxlpmlfklovrden <= '0';
      s_gth_rx_init_arr(i*4+j).RXDFELFOVRDEN   <= '0';
      s_gth_rx_init_arr(i*4+j).RXLPMHFOVRDEN   <= '0';

      --------------------------------------------------------------------------
      gt_cdrlock_timeout : process(clk_stable_i)
      begin
        if rising_edge(clk_stable_i) then
          if(gth_gt_rxreset_i(i*4+j) = '1') then
            s_gth_rx_cdrlocked(i*4+j)       <= '0';
            s_gth_rx_cdrlock_counter(i*4+j) <= 0;
          elsif (s_gth_rx_cdrlock_counter(i*4+j) = C_WAIT_TIME_CDRLOCK) then
            s_gth_rx_cdrlocked(i*4+j)       <= '1';
            s_gth_rx_cdrlock_counter(i*4+j) <= s_gth_rx_cdrlock_counter(i*4+j);
          else
            s_gth_rx_cdrlock_counter(i*4+j) <= s_gth_rx_cdrlock_counter(i*4+j) + 1;
          end if;
        end if;
      end process;

      s_gth_recclk_stable(i*4+j) <= s_gth_rx_cdrlocked(i*4+j);

      --------------------------- TX Buffer Bypass Logic --------------------
      -- The TX SYNC Module drives the ports needed to Bypass the TX Buffer.
      -- Include the TX SYNC module in your own design if TX Buffer is bypassed.

      --Manual
      i_gth_single_tx_manual_phase_align : entity work.gth_single_TX_MANUAL_PHASE_ALIGN
        generic map
        (
          NUMBER_OF_LANES => 1,
          MASTER_LANE_ID  => 0
          )
        port map
        (
          STABLE_CLOCK         => clk_stable_i,
          RESET_PHALIGNMENT    => s_gth_tx_rst_phalignment(i*4+j),  --TODO
          RUN_PHALIGNMENT      => s_gth_tx_run_phalignment(i*4+j),  --TODO
          PHASE_ALIGNMENT_DONE => s_gth_tx_run_phalignment_done(i*4+j),
          TXDLYSRESET(0)       => s_gth_tx_init_arr(i*4+j).TXDLYSRESET,
          TXDLYSRESETDONE(0)   => s_gth_tx_status_arr(i*4+j).TXDLYSRESETDONE,
          TXPHINIT(0)          => s_gth_tx_init_arr(i*4+j).TXPHINIT,
          TXPHINITDONE(0)      => s_gth_tx_status_arr(i*4+j).TXPHINITDONE,
          TXPHALIGN(0)         => s_gth_tx_init_arr(i*4+j).TXPHALIGN,
          TXPHALIGNDONE(0)     => s_gth_tx_status_arr(i*4+j).TXPHALIGNDONE,
          TXDLYEN(0)           => s_gth_tx_init_arr(i*4+j).TXDLYEN
          );
      s_gth_tx_init_arr(i*4+j).TXPHALIGNEN  <= '1';
      s_gth_tx_init_arr(i*4+j).TXPHDLYRESET <= '0';

      i_rx_auto_phase_align : entity work.gth_single_AUTO_PHASE_ALIGN
        port map (
          STABLE_CLOCK         => clk_stable_i,
          RUN_PHALIGNMENT      => s_gth_rx_run_phalignment(i*4+j),
          PHASE_ALIGNMENT_DONE => s_gth_rx_run_phalignment_done(i*4+j),
          PHALIGNDONE          => s_gth_rx_status_arr(i*4+j).RXSYNCDONE,
          DLYSRESET            => s_gth_rx_init_arr(i*4+j).RXDLYSRESET,
          DLYSRESETDONE        => s_gth_rx_status_arr(i*4+j).RXDLYSRESETDONE,
          RECCLKSTABLE         => s_gth_recclk_stable(i*4+j)
          );

      s_gth_rx_init_arr(i*4+j).RXCDRHOLD    <= '0';
      s_gth_rx_init_arr(i*4+j).RXPHDLYRESET <= '0';
      s_gth_rx_init_arr(i*4+j).RXPHALIGNEN  <= '0';
      s_gth_rx_init_arr(i*4+j).RXDLYEN      <= '0';
      s_gth_rx_init_arr(i*4+j).RXPHALIGN    <= '0';
      s_gth_rx_init_arr(i*4+j).RXSYNCMODE   <= '1';
      s_gth_rx_init_arr(i*4+j).RXSYNCIN     <= '0';
      s_gth_rx_init_arr(i*4+j).RXSYNCALLIN  <= s_gth_rx_status_arr(i*4+j).RXPHALIGNDONE;


    end generate;
  end generate;

end gth_wrapper_arch;
--============================================================================
--                                                            Architecture end
--============================================================================
